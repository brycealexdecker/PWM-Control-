** Profile: "SCHEMATIC1-TLV3231"  [ C:\Pspice Models\TLV3231\TLV3231-PSpice\TLV3231-PSpiceFiles\SCHEMATIC1\TLV3231.sim ] 

** Creating circuit file "TLV3231.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../tlv3231.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data-Silent\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:

*Analysis directives: 
.TRAN  0 30u 0 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
